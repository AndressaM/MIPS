module register_file( logic input A1[4:0], A2[4:0],A3[4:0] ,clk , logic output RD1,RD2);
	
endmodule