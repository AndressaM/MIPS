module main_controler(input logic [5:0]opcode ,
							output logic MentoReg,RegDst,IorD,
							PCSrc, output logic[1:0]ALUSrcB,ALUSrcA,IRWrite,
							MenWrite,PCWrite,Branch,RegWrite, output logic[1:0]ALUOp);
endmodule